library ieee;
use ieee.std_logic_1164.all;

entity COMPARADOR_10_BITS is
   port (A,B : in  std_logic_VECTOR(9 downto 0);
         QS : out std_logic); -- MAIOR OU IGUAL SERÁ O SINAL DE SAIDA
end COMPARADOR_10_BITS;

architecture CKT of COMPARADOR_10_BITS is

signal IGUAL : std_logic;
SIGNAL IGUAL9,IGUAL8,IGUAL7,IGUAL6,IGUAL5,IGUAL4,IGUAL3,IGUAL2,IGUAL1,IGUAL0 : std_logic;
SIGNAL IGUAL_8_9,IGUAL_7_9,IGUAL_6_9,IGUAL_5_9,IGUAL_4_9,IGUAL_3_9,IGUAL_2_9,IGUAL_1_9 : std_logic;
signal SAIDA1 : std_logic;

begin
IGUAL9 <= NOT(A(9) OR B(9));
IGUAL8 <= NOT(A(8) OR B(8));
IGUAL7 <= NOT(A(7) OR B(7));
IGUAL6 <= NOT(A(6) OR B(6));
IGUAL5 <= NOT(A(5) OR B(5));
IGUAL4 <= NOT(A(4) OR B(4));
IGUAL3 <= NOT(A(3) OR B(3));
IGUAL2 <= NOT(A(2) OR B(2));
IGUAL1 <= NOT(A(1) OR B(1));
IGUAL0 <= NOT(A(0) OR B(0));
IGUAL	 <= (IGUAL9 AND IGUAL8 AND IGUAL7 AND IGUAL6 AND IGUAL5 AND IGUAL4 AND IGUAL3 AND IGUAL2 AND IGUAL1 AND IGUAL0);
		
IGUAL_8_9	<= IGUAL9 AND IGUAL8;
IGUAL_7_9	<= IGUAL9 AND IGUAL8 AND IGUAL7;
IGUAL_6_9	<= IGUAL9 AND IGUAL8 AND IGUAL7 AND IGUAL6;
IGUAL_5_9	<= IGUAL9 AND IGUAL8 AND IGUAL7 AND IGUAL6 AND IGUAL5;
IGUAL_4_9	<= IGUAL9 AND IGUAL8 AND IGUAL7 AND IGUAL6 AND IGUAL5 AND IGUAL4;
IGUAL_3_9	<= IGUAL9 AND IGUAL8 AND IGUAL7 AND IGUAL6 AND IGUAL5 AND IGUAL4 AND IGUAL3;
IGUAL_2_9	<= IGUAL9 AND IGUAL8 AND IGUAL7 AND IGUAL6 AND IGUAL5 AND IGUAL4 AND IGUAL3 AND IGUAL2;
IGUAL_1_9	<= IGUAL9 AND IGUAL8 AND IGUAL7 AND IGUAL6 AND IGUAL5 AND IGUAL4 AND IGUAL3 AND IGUAL2 AND IGUAL1;


   
SAIDA1 <=  (A(9) AND (NOT B(9))) OR (IGUAL9 AND A(8) AND (NOT B(8))) OR (IGUAL_8_9 AND A(7) AND (NOT  B(7))) OR (IGUAL_7_9 AND A(6) AND (NOT B(6))) OR (IGUAL_6_9 AND A(5) AND (NOT B(5))) OR (IGUAL_5_9 AND A(4) AND (NOT B(4))) OR (IGUAL_4_9 AND A(3) AND (NOT B(3))) OR (IGUAL_3_9 AND A(2) AND (NOT B(2))) OR (IGUAL_2_9 AND A(1) AND (NOT B(1))) OR (IGUAL_1_9 AND A(0) AND (NOT B(0))); 

QS <= SAIDA1 OR IGUAL;
	
	
end CKT;