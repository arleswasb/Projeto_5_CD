library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity REGISTRADOR_10_BITS is
   Port (clk, clr, set : in STD_LOGIC;
		E :  in STD_LOGIC_VECTOR(9 downto 0);
         	S : out STD_LOGIC_VECTOR(9 downto 0));
end REGISTRADOR_10_BITS;

architecture ckt of REGISTRADOR_10_BITS is

	component ffd is
		port (ck, clr, set, d : in  std_logic;
								  q : out std_logic);
	end component;

	

	begin
	
		FF9:ffd port map (clk,clr,set,E(9),S(9));
		FF8:ffd port map (clk,clr,set,E(8),S(8));
		FF7:ffd port map (clk,clr,set,E(7),S(7));
		FF6:ffd port map (clk,clr,set,E(6),S(6));
		FF5:ffd port map (clk,clr,set,E(5),S(5));
		FF4:ffd port map (clk,clr,set,E(4),S(4));
		FF3:ffd port map (clk,clr,set,E(3),S(3));
		FF2:ffd port map (clk,clr,set,E(2),S(2));
		FF1:ffd port map (clk,clr,set,E(1),S(1));
		FF0:ffd port map (clk,clr,set,E(0),S(0));


end ckt;